package apb_pkg;
event e1;
`include "/home/dvft0904/apb_sv_project/env/transaction.sv"
`include "/home/dvft0904/apb_sv_project/env/generator.sv"
`include "/home/dvft0904/apb_sv_project/env/driver.sv"
`include "/home/dvft0904/apb_sv_project/env/monitor.sv"
`include "/home/dvft0904/apb_sv_project/env/predictor.sv"
`include "/home/dvft0904/apb_sv_project/env/scoreboard.sv"
`include "/home/dvft0904/apb_sv_project/env/environment.sv"
`include "/home/dvft0904/apb_sv_project/test/test.sv"
endpackage





